module top_810026173_826291639_946996917_1246901
//module top_810222780_826291639_829556405_4392126
//module top_809698492_826291639_762447541_4392120
( n14 , n17 , n19 , n26 , n33 , n36 , n44 , n46 , n49 , 
n55 , n56 , n66 , n67 , n69 , n74 , n106 , n126 , n135 , n145 , 
n155 , n156 , n171 , n174 , n181 , n183 , n208 , n213 , n216 , n218 , 
n223 , n231 , n238 , n247 , n266 , n270 , n276 , n277 , n290 , n292 , 
n299 , n303 , n317 , n329 , n347 , n353 , n372 , n378 , n379 , n387 , 
n391 , n401 , n402 , n414 , n416 , n423 , n424 , n426 , n429 , n432 , 
n433 , n444 , n452 , n457 , n460 , n469 , n472 , n476 , n482 , n488 , 
n493 , n498 , n510 , n517 , n522 , n532 , n534 , n541 , n547 , n549 , 
n555 , n557 , n559 , n569 , n573 , n585 , n588 , n599 , n600 , n607 , 
n627 , n638 , n643 , n646 , n647 , n648 , n649 , n653 , n655 , n665 , 
n675 , n682 , n683 , n684 , n693 , n695 , n699 , n712 , n715 , n724 , 
n725 , n729 , n731 , n738 , n747 , n748 , n759 , n761 , n770 , n773 , 
n788 , n790 , n792 , n801 , n813 , n823 , n824 , n836 , n839 , n846 , 
n858 , n862 , n865 , n867 , n870 , n882 , n883 , n888 , n891 , n892 , 
n902 , n905 , n906 , n912 , n927 , n931 , n935 , n942 , n944 , n952 , 
n953 , n961 , n968 , n974 , n979 , n980 , n989 , n991 , n1000 , n1005 , 
n1012 , n1015 , n1016 , n1025 , n1030 , n1062 , n1067 , n1068 , n1103 , n1113 , 
n1119 , n1135 , n1138 , n1140 , n1142 , n1145 , n1149 , n1161 , n1162 , n1172 , 
n1175 , n1183 , n1191 , n1194 , n1199 , n1201 , n1202 , n1222 , n1234 , n1235 , 
n1237 , n1249 , n1255 , n1260 , n1263 , n1277 , n1278 , n1283 , n1296 , n1305 , 
n1315 , n1321 , n1330 , n1332 , n1338 , n1340 , n1341 , n1347 , n1348 , n1349 , 
n1351 , n1363 , n1369 , n1381 , n1383 , n1385 , n1393 , n1399 , n1407 , n1422 , 
n1425 , n1426 , n1435 , n1440 , n1453 , n1457 , n1460 , n1461 , n1463 , n1470 , 
n1481 , n1495 , n1498 , n1501 , n1502 , n1507 , n1525 , n1527 , n1530 , n1535 , 
n1537 , n1544 , n1556 , n1595 , n1597 , n1600 , n1601 , n1613 , n1622 , n1629 , 
n1633 , n1635 , n1642 , n1643 , n1654 , n1657 , n1660 , n1675 , n1677 , n1678 , 
n1683 , n1686 , n1688 , n1690 , n1707 , n1721 , n1727 , n1729 , n1731 , n1737 , 
n1743 , n1746 , n1747 , n1757 , n1763 , n1764 );
    input n14 , n17 , n26 , n36 , n46 , n49 , n66 , n69 , n155 , 
n171 , n183 , n213 , n223 , n247 , n266 , n277 , n303 , n329 , n347 , 
n353 , n379 , n391 , n402 , n414 , n424 , n433 , n444 , n469 , n472 , 
n498 , n555 , n557 , n585 , n600 , n607 , n649 , n653 , n655 , n675 , 
n682 , n684 , n693 , n695 , n729 , n738 , n747 , n761 , n788 , n801 , 
n839 , n862 , n870 , n882 , n906 , n927 , n931 , n952 , n953 , n961 , 
n968 , n1000 , n1062 , n1140 , n1145 , n1172 , n1222 , n1263 , n1296 , n1321 , 
n1332 , n1341 , n1351 , n1363 , n1381 , n1422 , n1435 , n1461 , n1501 , n1527 , 
n1530 , n1537 , n1544 , n1597 , n1622 , n1642 , n1643 , n1678 , n1707 , n1743 , 
n1747 , n1757 , n1763 , n1764 ;
    output n19 , n33 , n44 , n55 , n56 , n67 , n74 , n106 , n126 , 
n135 , n145 , n156 , n174 , n181 , n208 , n216 , n218 , n231 , n238 , 
n270 , n276 , n290 , n292 , n299 , n317 , n372 , n378 , n387 , n401 , 
n416 , n423 , n426 , n429 , n432 , n452 , n457 , n460 , n476 , n482 , 
n488 , n493 , n510 , n517 , n522 , n532 , n534 , n541 , n547 , n549 , 
n559 , n569 , n573 , n588 , n599 , n627 , n638 , n643 , n646 , n647 , 
n648 , n665 , n683 , n699 , n712 , n715 , n724 , n725 , n731 , n748 , 
n759 , n770 , n773 , n790 , n792 , n813 , n823 , n824 , n836 , n846 , 
n858 , n865 , n867 , n883 , n888 , n891 , n892 , n902 , n905 , n912 , 
n935 , n942 , n944 , n974 , n979 , n980 , n989 , n991 , n1005 , n1012 , 
n1015 , n1016 , n1025 , n1030 , n1067 , n1068 , n1103 , n1113 , n1119 , n1135 , 
n1138 , n1142 , n1149 , n1161 , n1162 , n1175 , n1183 , n1191 , n1194 , n1199 , 
n1201 , n1202 , n1234 , n1235 , n1237 , n1249 , n1255 , n1260 , n1277 , n1278 , 
n1283 , n1305 , n1315 , n1330 , n1338 , n1340 , n1347 , n1348 , n1349 , n1369 , 
n1383 , n1385 , n1393 , n1399 , n1407 , n1425 , n1426 , n1440 , n1453 , n1457 , 
n1460 , n1463 , n1470 , n1481 , n1495 , n1498 , n1502 , n1507 , n1525 , n1535 , 
n1556 , n1595 , n1600 , n1601 , n1613 , n1629 , n1633 , n1635 , n1654 , n1657 , 
n1660 , n1675 , n1677 , n1683 , n1686 , n1688 , n1690 , n1721 , n1727 , n1729 , 
n1731 , n1737 , n1746 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n11 , n12 , n13 , n15 , n16 , n18 , n20 , n21 , 
n22 , n23 , n24 , n25 , n27 , n28 , n29 , n30 , n31 , n32 , 
n34 , n35 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n45 , 
n47 , n48 , n50 , n51 , n52 , n53 , n54 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n68 , n70 , n71 , n72 , 
n73 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , 
n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , 
n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , 
n104 , n105 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , 
n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , 
n125 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n136 , 
n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n146 , n147 , 
n148 , n149 , n150 , n151 , n152 , n153 , n154 , n157 , n158 , n159 , 
n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
n170 , n172 , n173 , n175 , n176 , n177 , n178 , n179 , n180 , n182 , 
n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , 
n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , 
n204 , n205 , n206 , n207 , n209 , n210 , n211 , n212 , n214 , n215 , 
n217 , n219 , n220 , n221 , n222 , n224 , n225 , n226 , n227 , n228 , 
n229 , n230 , n232 , n233 , n234 , n235 , n236 , n237 , n239 , n240 , 
n241 , n242 , n243 , n244 , n245 , n246 , n248 , n249 , n250 , n251 , 
n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , 
n262 , n263 , n264 , n265 , n267 , n268 , n269 , n271 , n272 , n273 , 
n274 , n275 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , 
n286 , n287 , n288 , n289 , n291 , n293 , n294 , n295 , n296 , n297 , 
n298 , n300 , n301 , n302 , n304 , n305 , n306 , n307 , n308 , n309 , 
n310 , n311 , n312 , n313 , n314 , n315 , n316 , n318 , n319 , n320 , 
n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n330 , n331 , 
n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , 
n342 , n343 , n344 , n345 , n346 , n348 , n349 , n350 , n351 , n352 , 
n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , 
n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n373 , n374 , 
n375 , n376 , n377 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
n388 , n389 , n390 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , 
n399 , n400 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
n411 , n412 , n413 , n415 , n417 , n418 , n419 , n420 , n421 , n422 , 
n425 , n427 , n428 , n430 , n431 , n434 , n435 , n436 , n437 , n438 , 
n439 , n440 , n441 , n442 , n443 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n453 , n454 , n455 , n456 , n458 , n459 , n461 , n462 , 
n463 , n464 , n465 , n466 , n467 , n468 , n470 , n471 , n473 , n474 , 
n475 , n477 , n478 , n479 , n480 , n481 , n483 , n484 , n485 , n486 , 
n487 , n489 , n490 , n491 , n492 , n494 , n495 , n496 , n497 , n499 , 
n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n511 , n512 , n513 , n514 , n515 , n516 , n518 , n519 , n520 , n521 , 
n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n533 , 
n535 , n536 , n537 , n538 , n539 , n540 , n542 , n543 , n544 , n545 , 
n546 , n548 , n550 , n551 , n552 , n553 , n554 , n556 , n558 , n560 , 
n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n570 , n571 , 
n572 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , 
n583 , n584 , n586 , n587 , n589 , n590 , n591 , n592 , n593 , n594 , 
n595 , n596 , n597 , n598 , n601 , n602 , n603 , n604 , n605 , n606 , 
n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , 
n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n628 , 
n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n639 , 
n640 , n641 , n642 , n644 , n645 , n650 , n651 , n652 , n654 , n656 , 
n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n666 , n667 , 
n668 , n669 , n670 , n671 , n672 , n673 , n674 , n676 , n677 , n678 , 
n679 , n680 , n681 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , 
n692 , n694 , n696 , n697 , n698 , n700 , n701 , n702 , n703 , n704 , 
n705 , n706 , n707 , n708 , n709 , n710 , n711 , n713 , n714 , n716 , 
n717 , n718 , n719 , n720 , n721 , n722 , n723 , n726 , n727 , n728 , 
n730 , n732 , n733 , n734 , n735 , n736 , n737 , n739 , n740 , n741 , 
n742 , n743 , n744 , n745 , n746 , n749 , n750 , n751 , n752 , n753 , 
n754 , n755 , n756 , n757 , n758 , n760 , n762 , n763 , n764 , n765 , 
n766 , n767 , n768 , n769 , n771 , n772 , n774 , n775 , n776 , n777 , 
n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , 
n789 , n791 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , 
n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , 
n812 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , 
n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , 
n835 , n837 , n838 , n840 , n841 , n842 , n843 , n844 , n845 , n847 , 
n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , 
n859 , n860 , n861 , n863 , n864 , n866 , n868 , n869 , n871 , n872 , 
n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n884 , 
n885 , n886 , n887 , n889 , n890 , n893 , n894 , n895 , n896 , n897 , 
n898 , n899 , n900 , n901 , n903 , n904 , n907 , n908 , n909 , n910 , 
n911 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , 
n922 , n923 , n924 , n925 , n926 , n928 , n929 , n930 , n932 , n933 , 
n934 , n936 , n937 , n938 , n939 , n940 , n941 , n943 , n945 , n946 , 
n947 , n948 , n949 , n950 , n951 , n954 , n955 , n956 , n957 , n958 , 
n959 , n960 , n962 , n963 , n964 , n965 , n966 , n967 , n969 , n970 , 
n971 , n972 , n973 , n975 , n976 , n977 , n978 , n981 , n982 , n983 , 
n984 , n985 , n986 , n987 , n988 , n990 , n992 , n993 , n994 , n995 , 
n996 , n997 , n998 , n999 , n1001 , n1002 , n1003 , n1004 , n1006 , n1007 , 
n1008 , n1009 , n1010 , n1011 , n1013 , n1014 , n1017 , n1018 , n1019 , n1020 , 
n1021 , n1022 , n1023 , n1024 , n1026 , n1027 , n1028 , n1029 , n1031 , n1032 , 
n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , 
n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , 
n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1063 , 
n1064 , n1065 , n1066 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , 
n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , 
n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , 
n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1104 , n1105 , n1106 , 
n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1114 , n1115 , n1116 , n1117 , 
n1118 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , 
n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1136 , n1137 , n1139 , n1141 , 
n1143 , n1144 , n1146 , n1147 , n1148 , n1150 , n1151 , n1152 , n1153 , n1154 , 
n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1163 , n1164 , n1165 , n1166 , 
n1167 , n1168 , n1169 , n1170 , n1171 , n1173 , n1174 , n1176 , n1177 , n1178 , 
n1179 , n1180 , n1181 , n1182 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
n1190 , n1192 , n1193 , n1195 , n1196 , n1197 , n1198 , n1200 , n1203 , n1204 , 
n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , 
n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1223 , n1224 , n1225 , 
n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1236 , n1238 , 
n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , 
n1250 , n1251 , n1252 , n1253 , n1254 , n1256 , n1257 , n1258 , n1259 , n1261 , 
n1262 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , 
n1273 , n1274 , n1275 , n1276 , n1279 , n1280 , n1281 , n1282 , n1284 , n1285 , 
n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , 
n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1306 , n1307 , 
n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1316 , n1317 , n1318 , 
n1319 , n1320 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1331 , n1333 , n1334 , n1335 , n1336 , n1337 , n1339 , n1342 , n1343 , n1344 , 
n1345 , n1346 , n1350 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , 
n1359 , n1360 , n1361 , n1362 , n1364 , n1365 , n1366 , n1367 , n1368 , n1370 , 
n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
n1382 , n1384 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1394 , 
n1395 , n1396 , n1397 , n1398 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , 
n1406 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , 
n1417 , n1418 , n1419 , n1420 , n1421 , n1423 , n1424 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1436 , n1437 , n1438 , n1439 , n1441 , 
n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , 
n1452 , n1454 , n1455 , n1456 , n1458 , n1459 , n1462 , n1464 , n1465 , n1466 , 
n1467 , n1468 , n1469 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , 
n1478 , n1479 , n1480 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , 
n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1496 , n1497 , n1499 , n1500 , 
n1503 , n1504 , n1505 , n1506 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , 
n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , 
n1524 , n1526 , n1528 , n1529 , n1531 , n1532 , n1533 , n1534 , n1536 , n1538 , 
n1539 , n1540 , n1541 , n1542 , n1543 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1557 , n1558 , n1559 , n1560 , 
n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
n1591 , n1592 , n1593 , n1594 , n1596 , n1598 , n1599 , n1602 , n1603 , n1604 , 
n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1614 , n1615 , 
n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1623 , n1624 , n1625 , n1626 , 
n1627 , n1628 , n1630 , n1631 , n1632 , n1634 , n1636 , n1637 , n1638 , n1639 , 
n1640 , n1641 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , 
n1652 , n1653 , n1655 , n1656 , n1658 , n1659 , n1661 , n1662 , n1663 , n1664 , 
n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , 
n1676 , n1679 , n1680 , n1681 , n1682 , n1684 , n1685 , n1687 , n1689 , n1691 , 
n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , 
n1702 , n1703 , n1704 , n1705 , n1706 , n1708 , n1709 , n1710 , n1711 , n1712 , 
n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1722 , n1723 , 
n1724 , n1725 , n1726 , n1728 , n1730 , n1732 , n1733 , n1734 , n1735 , n1736 , 
n1738 , n1739 , n1740 , n1741 , n1742 , n1744 , n1745 , n1748 , n1749 , n1750 , 
n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1758 , n1759 , n1760 , n1761 , 
n1762 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 ;
    or g0 ( n1251 , n235 , n1266 );
    not g1 ( n1565 , n527 );
    not g2 ( n1312 , n1653 );
    or g3 ( n1414 , n1090 , n673 );
    xnor g4 ( n1352 , n298 , n1568 );
    xnor g5 ( n599 , n416 , n1403 );
    or g6 ( n1037 , n188 , n554 );
    nor g7 ( n540 , n654 , n986 );
    or g8 ( n1181 , n1582 , n72 );
    or g9 ( n473 , n562 , n1653 );
    not g10 ( n1146 , n911 );
    xnor g11 ( n1432 , n265 , n953 );
    and g12 ( n188 , n952 , n329 );
    xnor g13 ( n229 , n283 , n557 );
    and g14 ( n13 , n1085 , n1290 );
    and g15 ( n1272 , n1312 , n214 );
    not g16 ( n1716 , n390 );
    and g17 ( n361 , n1429 , n1126 );
    xnor g18 ( n1523 , n1390 , n1645 );
    and g19 ( n702 , n1750 , n582 );
    nor g20 ( n1368 , n1343 , n816 );
    nor g21 ( n662 , n1371 , n1169 );
    xnor g22 ( n1015 , n960 , n458 );
    or g23 ( n1156 , n874 , n193 );
    or g24 ( n696 , n1263 , n1444 );
    or g25 ( n1596 , n1316 , n316 );
    and g26 ( n827 , n1255 , n1155 );
    or g27 ( n1079 , n441 , n264 );
    xnor g28 ( n1502 , n255 , n727 );
    and g29 ( n1725 , n898 , n1171 );
    and g30 ( n1318 , n1692 , n589 );
    nor g31 ( n1384 , n1174 , n48 );
    nor g32 ( n744 , n257 , n552 );
    and g33 ( n1697 , n101 , n283 );
    or g34 ( n308 , n1170 , n392 );
    or g35 ( n78 , n326 , n1680 );
    not g36 ( n1634 , n1282 );
    xnor g37 ( n1391 , n128 , n92 );
    xnor g38 ( n1003 , n1607 , n1764 );
    xnor g39 ( n20 , n1671 , n305 );
    and g40 ( n1664 , n473 , n1404 );
    not g41 ( n1410 , n722 );
    xnor g42 ( n1155 , n962 , n259 );
    or g43 ( n88 , n1527 , n46 );
    and g44 ( n228 , n1409 , n1099 );
    or g45 ( n458 , n96 , n698 );
    or g46 ( n1499 , n1642 , n1232 );
    xnor g47 ( n1234 , n1458 , n569 );
    or g48 ( n35 , n543 , n706 );
    xnor g49 ( n726 , n816 , n1579 );
    and g50 ( n819 , n1622 , n1346 );
    and g51 ( n12 , n922 , n1508 );
    or g52 ( n485 , n1057 , n463 );
    not g53 ( n704 , n1037 );
    not g54 ( n1770 , n1104 );
    and g55 ( n434 , n202 , n1276 );
    and g56 ( n63 , n503 , n1547 );
    xnor g57 ( n846 , n604 , n286 );
    and g58 ( n1602 , n227 , n367 );
    and g59 ( n580 , n1727 , n1663 );
    xnor g60 ( n1046 , n1643 , n1707 );
    not g61 ( n1773 , n1007 );
    nor g62 ( n1722 , n164 , n347 );
    and g63 ( n1702 , n1461 , n1381 );
    xnor g64 ( n665 , n831 , n1698 );
    or g65 ( n1756 , n1734 , n1639 );
    not g66 ( n1174 , n123 );
    not g67 ( n843 , n133 );
    not g68 ( n529 , n119 );
    not g69 ( n398 , n936 );
    xnor g70 ( n902 , n1099 , n1359 );
    nor g71 ( n925 , n1768 , n1167 );
    xnor g72 ( n1005 , n125 , n103 );
    not g73 ( n1647 , n331 );
    or g74 ( n146 , n1381 , n1116 );
    nor g75 ( n1715 , n555 , n1014 );
    not g76 ( n125 , n550 );
    xnor g77 ( n1609 , n1254 , n243 );
    or g78 ( n192 , n1329 , n266 );
    xnor g79 ( n1398 , n5 , n260 );
    xnor g80 ( n428 , n16 , n254 );
    xnor g81 ( n1730 , n815 , n1357 );
    xnor g82 ( n1284 , n1204 , n112 );
    not g83 ( n1322 , n203 );
    not g84 ( n584 , n362 );
    and g85 ( n1614 , n1337 , n131 );
    and g86 ( n1739 , n1658 , n179 );
    not g87 ( n371 , n682 );
    nor g88 ( n42 , n1442 , n994 );
    not g89 ( n1366 , n1363 );
    nor g90 ( n947 , n195 , n565 );
    or g91 ( n367 , n1381 , n601 );
    not g92 ( n73 , n1578 );
    and g93 ( n1243 , n1511 , n1767 );
    and g94 ( n1173 , n1473 , n1769 );
    xnor g95 ( n387 , n1271 , n1425 );
    or g96 ( n834 , n789 , n249 );
    not g97 ( n474 , n954 );
    not g98 ( n1018 , n111 );
    and g99 ( n1456 , n382 , n474 );
    nor g100 ( n443 , n46 , n805 );
    or g101 ( n1327 , n1381 , n309 );
    xnor g102 ( n1762 , n1146 , n497 );
    and g103 ( n639 , n1566 , n1771 );
    nor g104 ( n1090 , n1442 , n1335 );
    nor g105 ( n590 , n1643 , n1709 );
    not g106 ( n157 , n953 );
    xnor g107 ( n1106 , n268 , n486 );
    or g108 ( n901 , n1626 , n1164 );
    xnor g109 ( n1688 , n1168 , n898 );
    or g110 ( n470 , n605 , n548 );
    and g111 ( n1147 , n568 , n1076 );
    not g112 ( n177 , n379 );
    and g113 ( n535 , n472 , n99 );
    and g114 ( n921 , n332 , n1055 );
    or g115 ( n258 , n1543 , n233 );
    nor g116 ( n77 , n1469 , n558 );
    and g117 ( n338 , n1100 , n826 );
    or g118 ( n1317 , n1219 , n312 );
    not g119 ( n312 , n1280 );
    or g120 ( n767 , n820 , n1167 );
    or g121 ( n924 , n895 , n596 );
    or g122 ( n911 , n1323 , n640 );
    or g123 ( n158 , n1532 , n1472 );
    xnor g124 ( n857 , n99 , n1743 );
    and g125 ( n108 , n1684 , n39 );
    and g126 ( n539 , n1112 , n1048 );
    not g127 ( n715 , n1408 );
    xnor g128 ( n368 , n1443 , n213 );
    xnor g129 ( n55 , n626 , n898 );
    not g130 ( n408 , n275 );
    or g131 ( n1211 , n40 , n75 );
    nor g132 ( n1388 , n1259 , n593 );
    and g133 ( n1486 , n1678 , n1381 );
    nor g134 ( n971 , n1065 , n1598 );
    not g135 ( n1268 , n1420 );
    not g136 ( n536 , n810 );
    or g137 ( n1606 , n57 , n1685 );
    buf g138 ( n174 , n488 );
    not g139 ( n708 , n449 );
    xnor g140 ( n582 , n1709 , n1474 );
    or g141 ( n1259 , n1310 , n1590 );
    or g142 ( n1517 , n102 , n191 );
    or g143 ( n129 , n562 , n73 );
    and g144 ( n370 , n1121 , n1367 );
    nor g145 ( n160 , n952 , n197 );
    xnor g146 ( n1353 , n275 , n600 );
    and g147 ( n1210 , n1261 , n611 );
    or g148 ( n212 , n175 , n1374 );
    or g149 ( n278 , n947 , n1567 );
    and g150 ( n1719 , n827 , n1244 );
    nor g151 ( n1621 , n876 , n570 );
    not g152 ( n676 , n495 );
    or g153 ( n1242 , n1497 , n1061 );
    and g154 ( n749 , n391 , n536 );
    nor g155 ( n1245 , n1642 , n1617 );
    or g156 ( n1367 , n10 , n12 );
    xnor g157 ( n1407 , n673 , n1733 );
    xnor g158 ( n1302 , n1057 , n1169 );
    not g159 ( n1320 , n753 );
    and g160 ( n90 , n295 , n1215 );
    not g161 ( n1700 , n1592 );
    not g162 ( n809 , n839 );
    not g163 ( n669 , n70 );
    and g164 ( n1586 , n226 , n386 );
    or g165 ( n946 , n1532 , n296 );
    not g166 ( n1082 , n1115 );
    xnor g167 ( n849 , n633 , n303 );
    not g168 ( n1119 , n471 );
    and g169 ( n1449 , n1435 , n1532 );
    not g170 ( n735 , n1448 );
    not g171 ( n820 , n247 );
    not g172 ( n1316 , n1381 );
    or g173 ( n570 , n667 , n166 );
    and g174 ( n938 , n1435 , n1167 );
    xor g175 ( n1641 , n1274 , n247 );
    xnor g176 ( n376 , n1512 , n1581 );
    or g177 ( n863 , n164 , n1381 );
    not g178 ( n710 , n1571 );
    and g179 ( n1550 , n657 , n308 );
    or g180 ( n807 , n94 , n1405 );
    and g181 ( n1324 , n926 , n211 );
    not g182 ( n1749 , n288 );
    xnor g183 ( n170 , n1606 , n1222 );
    and g184 ( n1323 , n1381 , n1101 );
    and g185 ( n1054 , n1063 , n1414 );
    and g186 ( n374 , n1084 , n244 );
    or g187 ( n70 , n301 , n1506 );
    and g188 ( n45 , n978 , n924 );
    nor g189 ( n237 , n353 , n655 );
    nor g190 ( n534 , n923 , n660 );
    nor g191 ( n68 , n397 , n769 );
    and g192 ( n714 , n1044 , n995 );
    or g193 ( n1563 , n166 , n1353 );
    xnor g194 ( n1639 , n1120 , n437 );
    and g195 ( n169 , n360 , n998 );
    or g196 ( n124 , n262 , n361 );
    or g197 ( n1365 , n23 , n996 );
    not g198 ( n654 , n737 );
    not g199 ( n915 , n1456 );
    xnor g200 ( n648 , n511 , n1352 );
    and g201 ( n53 , n869 , n350 );
    not g202 ( n1637 , n1062 );
    not g203 ( n366 , n16 );
    xnor g204 ( n687 , n1607 , n1062 );
    xnor g205 ( n1463 , n28 , n139 );
    and g206 ( n1455 , n738 , n1485 );
    or g207 ( n246 , n366 , n137 );
    or g208 ( n932 , n579 , n354 );
    xnor g209 ( n76 , n1673 , n133 );
    nor g210 ( n148 , n863 , n1611 );
    not g211 ( n235 , n1527 );
    nor g212 ( n1292 , n1469 , n1111 );
    or g213 ( n541 , n829 , n527 );
    and g214 ( n22 , n413 , n764 );
    and g215 ( n122 , n1416 , n701 );
    and g216 ( n1539 , n720 , n185 );
    or g217 ( n873 , n711 , n908 );
    or g218 ( n487 , n343 , n1606 );
    nor g219 ( n121 , n223 , n1584 );
    not g220 ( n71 , n1224 );
    or g221 ( n1084 , n1287 , n1528 );
    or g222 ( n826 , n110 , n1594 );
    nor g223 ( n442 , n1217 , n679 );
    or g224 ( n325 , n1082 , n1639 );
    xnor g225 ( n1349 , n1239 , n1373 );
    not g226 ( n1385 , n614 );
    not g227 ( n659 , n787 );
    nor g228 ( n1053 , n253 , n1042 );
    xnor g229 ( n1280 , n326 , n93 );
    xnor g230 ( n522 , n323 , n352 );
    xnor g231 ( n1149 , n652 , n851 );
    not g232 ( n322 , n1480 );
    not g233 ( n561 , n112 );
    or g234 ( n1112 , n1568 , n298 );
    xnor g235 ( n1065 , n780 , n277 );
    or g236 ( n422 , n79 , n1627 );
    not g237 ( n96 , n1601 );
    and g238 ( n1182 , n1544 , n749 );
    and g239 ( n1477 , n806 , n1117 );
    nor g240 ( n903 , n952 , n265 );
    nor g241 ( n477 , n1597 , n266 );
    xnor g242 ( n1304 , n1300 , n271 );
    not g243 ( n742 , n1636 );
    and g244 ( n996 , n219 , n395 );
    or g245 ( n642 , n825 , n832 );
    or g246 ( n586 , n1316 , n269 );
    or g247 ( n1121 , n291 , n1089 );
    not g248 ( n382 , n1185 );
    or g249 ( n754 , n1604 , n234 );
    or g250 ( n1040 , n1422 , n696 );
    not g251 ( n764 , n1762 );
    xnor g252 ( n462 , n952 , n653 );
    xnor g253 ( n234 , n507 , n796 );
    not g254 ( n777 , n763 );
    xnor g255 ( n1676 , n1266 , n4 );
    and g256 ( n525 , n1386 , n631 );
    not g257 ( n825 , n1115 );
    or g258 ( n840 , n533 , n1662 );
    xnor g259 ( n1213 , n1154 , n862 );
    or g260 ( n1286 , n1344 , n704 );
    or g261 ( n810 , n1328 , n453 );
    not g262 ( n1685 , n1154 );
    not g263 ( n271 , n75 );
    or g264 ( n1279 , n1585 , n279 );
    xnor g265 ( n948 , n1604 , n1169 );
    and g266 ( n943 , n1694 , n1638 );
    not g267 ( n1342 , n797 );
    xnor g268 ( n748 , n1203 , n242 );
    not g269 ( n1503 , n246 );
    not g270 ( n1769 , n1519 );
    xnor g271 ( n890 , n1576 , n46 );
    or g272 ( n1511 , n490 , n281 );
    xnor g273 ( n1068 , n1391 , n1755 );
    or g274 ( n664 , n322 , n407 );
    xnor g275 ( n306 , n1575 , n736 );
    xnor g276 ( n1165 , n1602 , n390 );
    xnor g277 ( n759 , n30 , n1766 );
    xnor g278 ( n1475 , n73 , n200 );
    not g279 ( n1138 , n284 );
    not g280 ( n851 , n78 );
    xnor g281 ( n1201 , n1331 , n1714 );
    xnor g282 ( n951 , n1365 , n693 );
    and g283 ( n190 , n141 , n1038 );
    not g284 ( n869 , n721 );
    buf g285 ( n898 , n438 );
    nor g286 ( n47 , n1643 , n36 );
    xnor g287 ( n1199 , n644 , n215 );
    xnor g288 ( n51 , n1190 , n1708 );
    or g289 ( n611 , n853 , n1054 );
    xnor g290 ( n260 , n1618 , n1763 );
    not g291 ( n448 , n411 );
    and g292 ( n595 , n1652 , n60 );
    not g293 ( n889 , n856 );
    or g294 ( n1126 , n1510 , n415 );
    not g295 ( n200 , n1225 );
    or g296 ( n84 , n1316 , n618 );
    or g297 ( n481 , n272 , n1102 );
    nor g298 ( n321 , n447 , n516 );
    xnor g299 ( n305 , n1034 , n1643 );
    xnor g300 ( n1023 , n555 , n1172 );
    or g301 ( n597 , n164 , n574 );
    nor g302 ( n514 , n654 , n692 );
    or g303 ( n98 , n80 , n551 );
    nor g304 ( n551 , n563 , n1306 );
    or g305 ( n454 , n1479 , n576 );
    xnor g306 ( n208 , n994 , n117 );
    xnor g307 ( n1081 , n39 , n1684 );
    xnor g308 ( n1684 , n27 , n738 );
    xnor g309 ( n888 , n1567 , n1552 );
    and g310 ( n144 , n1073 , n934 );
    xnor g311 ( n44 , n1731 , n87 );
    nor g312 ( n484 , n1371 , n1555 );
    and g313 ( n1333 , n1259 , n436 );
    or g314 ( n173 , n1666 , n1710 );
    not g315 ( n916 , n819 );
    xnor g316 ( n65 , n1014 , n555 );
    or g317 ( n113 , n1532 , n1593 );
    not g318 ( n1184 , n1483 );
    not g319 ( n1558 , n1501 );
    not g320 ( n1665 , n718 );
    not g321 ( n0 , n1763 );
    nor g322 ( n1588 , n722 , n1717 );
    and g323 ( n1001 , n1394 , n1141 );
    or g324 ( n41 , n1195 , n75 );
    nor g325 ( n1047 , n1473 , n1769 );
    nor g326 ( n1509 , n1275 , n1751 );
    nor g327 ( n976 , n199 , n1531 );
    or g328 ( n546 , n1588 , n190 );
    or g329 ( n345 , n794 , n758 );
    xnor g330 ( n1030 , n1180 , n1326 );
    xnor g331 ( n900 , n1207 , n31 );
    and g332 ( n1216 , n578 , n1156 );
    xnor g333 ( n1560 , n720 , n1370 );
    or g334 ( n1459 , n1146 , n1004 );
    or g335 ( n1418 , n535 , n68 );
    not g336 ( n1070 , n489 );
    not g337 ( n523 , n1014 );
    or g338 ( n1694 , n509 , n1505 );
    xnor g339 ( n1582 , n1240 , n1332 );
    and g340 ( n50 , n969 , n1184 );
    and g341 ( n1289 , n222 , n1008 );
    xnor g342 ( n572 , n203 , n1579 );
    xnor g343 ( n731 , n63 , n1676 );
    xnor g344 ( n400 , n969 , n1483 );
    nor g345 ( n1295 , n584 , n1354 );
    xnor g346 ( n617 , n620 , n803 );
    and g347 ( n1116 , n206 , n597 );
    or g348 ( n456 , n1139 , n832 );
    not g349 ( n1029 , n1748 );
    xnor g350 ( n482 , n13 , n194 );
    xnor g351 ( n352 , n879 , n268 );
    and g352 ( n1620 , n171 , n1499 );
    not g353 ( n39 , n861 );
    or g354 ( n393 , n1000 , n1040 );
    xnor g355 ( n1729 , n998 , n1049 );
    xnor g356 ( n1230 , n1564 , n1544 );
    and g357 ( n497 , n1250 , n1534 );
    not g358 ( n395 , n1618 );
    and g359 ( n604 , n1400 , n267 );
    and g360 ( n1592 , n1034 , n1129 );
    xnor g361 ( n1064 , n24 , n781 );
    xnor g362 ( n449 , n412 , n1661 );
    xnor g363 ( n409 , n555 , n1140 );
    xnor g364 ( n1425 , n1673 , n1108 );
    and g365 ( n254 , n528 , n1433 );
    or g366 ( n1050 , n232 , n894 );
    not g367 ( n268 , n1284 );
    nor g368 ( n980 , n1084 , n1272 );
    xnor g369 ( n1690 , n118 , n610 );
    or g370 ( n1133 , n886 , n1137 );
    and g371 ( n1546 , n1317 , n431 );
    not g372 ( n9 , n832 );
    nor g373 ( n1220 , n741 , n1158 );
    and g374 ( n627 , n824 , n1271 );
    nor g375 ( n349 , n1208 , n104 );
    not g376 ( n1129 , n637 );
    not g377 ( n351 , n658 );
    nor g378 ( n496 , n121 , n1216 );
    not g379 ( n32 , n501 );
    not g380 ( n493 , n1078 );
    not g381 ( n241 , n393 );
    and g382 ( n1319 , n1124 , n1650 );
    not g383 ( n1013 , n994 );
    xnor g384 ( n1031 , n454 , n1432 );
    not g385 ( n1457 , n1609 );
    xnor g386 ( n1595 , n990 , n1348 );
    nor g387 ( n524 , n1513 , n402 );
    nor g388 ( n1467 , n478 , n475 );
    and g389 ( n973 , n1533 , n412 );
    not g390 ( n1346 , n987 );
    xnor g391 ( n1135 , n35 , n1333 );
    xnor g392 ( n33 , n639 , n273 );
    xnor g393 ( n1451 , n1082 , n351 );
    not g394 ( n1667 , n698 );
    not g395 ( n1576 , n163 );
    not g396 ( n802 , n695 );
    and g397 ( n153 , n34 , n1728 );
    nor g398 ( n287 , n855 , n1671 );
    xnor g399 ( n883 , n1165 , n1074 );
    not g400 ( n1099 , n1353 );
    and g401 ( n1334 , n1741 , n774 );
    and g402 ( n814 , n682 , n1371 );
    nor g403 ( n618 , n1620 , n283 );
    and g404 ( n1239 , n456 , n808 );
    not g405 ( n1115 , n123 );
    or g406 ( n830 , n1381 , n615 );
    not g407 ( n339 , n838 );
    and g408 ( n928 , n1568 , n298 );
    xnor g409 ( n1657 , n2 , n1138 );
    not g410 ( n530 , n607 );
    xnor g411 ( n452 , n1273 , n1523 );
    nor g412 ( n479 , n555 , n1172 );
    nor g413 ( n717 , n852 , n1052 );
    and g414 ( n249 , n957 , n1679 );
    or g415 ( n222 , n1723 , n1505 );
    or g416 ( n112 , n972 , n1018 );
    not g417 ( n641 , n54 );
    xnor g418 ( n786 , n353 , n655 );
    and g419 ( n1376 , n906 , n819 );
    xnor g420 ( n858 , n1491 , n500 );
    not g421 ( n1492 , n1444 );
    xnor g422 ( n1430 , n98 , n353 );
    nor g423 ( n750 , n1324 , n616 );
    nor g424 ( n1130 , n101 , n402 );
    or g425 ( n1100 , n359 , n1374 );
    nor g426 ( n1669 , n1322 , n228 );
    or g427 ( n189 , n101 , n335 );
    nor g428 ( n1476 , n1265 , n795 );
    xnor g429 ( n307 , n797 , n433 );
    and g430 ( n1720 , n1300 , n1581 );
    or g431 ( n1369 , n864 , n1333 );
    and g432 ( n1594 , n955 , n1454 );
    or g433 ( n1087 , n737 , n302 );
    xnor g434 ( n1552 , n435 , n195 );
    xnor g435 ( n1372 , n1217 , n379 );
    and g436 ( n316 , n723 , n1232 );
    nor g437 ( n811 , n585 , n402 );
    xnor g438 ( n1161 , n1141 , n828 );
    and g439 ( n451 , n505 , n933 );
    or g440 ( n528 , n1691 , n477 );
    xnor g441 ( n727 , n104 , n1480 );
    and g442 ( n1711 , n543 , n1224 );
    not g443 ( n1542 , n464 );
    xnor g444 ( n1077 , n197 , n472 );
    or g445 ( n204 , n1152 , n1327 );
    not g446 ( n293 , n696 );
    or g447 ( n1420 , n1051 , n775 );
    nor g448 ( n1699 , n66 , n1442 );
    and g449 ( n1528 , n91 , n144 );
    not g450 ( n1257 , n1190 );
    not g451 ( n871 , n1617 );
    or g452 ( n1378 , n240 , n620 );
    and g453 ( n824 , n1093 , n1724 );
    not g454 ( n511 , n122 );
    xnor g455 ( n194 , n825 , n48 );
    and g456 ( n1659 , n177 , n88 );
    not g457 ( n917 , n396 );
    not g458 ( n1445 , n1105 );
    nor g459 ( n1091 , n667 , n266 );
    and g460 ( n1608 , n223 , n1584 );
    not g461 ( n217 , n1474 );
    not g462 ( n1249 , n711 );
    and g463 ( n1011 , n1177 , n1110 );
    and g464 ( n673 , n833 , n1096 );
    or g465 ( n1709 , n1486 , n384 );
    or g466 ( n1580 , n177 , n879 );
    xnor g467 ( n818 , n1450 , n587 );
    or g468 ( n762 , n659 , n312 );
    and g469 ( n1331 , n1231 , n251 );
    xnor g470 ( n56 , n1143 , n172 );
    or g471 ( n1437 , n1607 , n440 );
    nor g472 ( n1488 , n1217 , n1280 );
    and g473 ( n757 , n1375 , n331 );
    xnor g474 ( n680 , n338 , n65 );
    nor g475 ( n1589 , n257 , n1725 );
    nor g476 ( n743 , n1461 , n402 );
    not g477 ( n1512 , n489 );
    or g478 ( n1765 , n486 , n268 );
    or g479 ( n1753 , n1695 , n209 );
    and g480 ( n100 , n1708 , n1257 );
    and g481 ( n678 , n1580 , n1738 );
    not g482 ( n83 , n849 );
    or g483 ( n1741 , n1415 , n658 );
    nor g484 ( n1308 , n624 , n1147 );
    or g485 ( n202 , n1300 , n72 );
    and g486 ( n1401 , n675 , n1214 );
    xnor g487 ( n432 , n233 , n773 );
    xnor g488 ( n711 , n1307 , n1397 );
    or g489 ( n336 , n413 , n764 );
    or g490 ( n131 , n1699 , n21 );
    nor g491 ( n1471 , n543 , n1224 );
    and g492 ( n209 , n1269 , n118 );
    not g493 ( n1673 , n1093 );
    xnor g494 ( n815 , n361 , n1021 );
    xnor g495 ( n460 , n1605 , n728 );
    xnor g496 ( n573 , n1625 , n948 );
    or g497 ( n1613 , n591 , n1658 );
    xnor g498 ( n274 , n447 , n1084 );
    and g499 ( n30 , n336 , n765 );
    nor g500 ( n583 , n1768 , n402 );
    xnor g501 ( n500 , n1581 , n1265 );
    and g502 ( n829 , n1721 , n406 );
    nor g503 ( n300 , n447 , n1312 );
    and g504 ( n548 , n860 , n1605 );
    xnor g505 ( n1473 , n1437 , n462 );
    or g506 ( n1496 , n504 , n676 );
    nor g507 ( n1759 , n953 , n265 );
    or g508 ( n227 , n1316 , n229 );
    not g509 ( n1223 , n960 );
    nor g510 ( n1392 , n1371 , n1645 );
    not g511 ( n291 , n555 );
    xnor g512 ( n935 , n1149 , n162 );
    not g513 ( n165 , n252 );
    or g514 ( n995 , n1043 , n1075 );
    not g515 ( n733 , n1499 );
    or g516 ( n616 , n164 , n355 );
    xnor g517 ( n1556 , n1426 , n96 );
    nor g518 ( n800 , n1217 , n268 );
    xnor g519 ( n1364 , n678 , n1166 );
    xnor g520 ( n273 , n509 , n1357 );
    or g521 ( n346 , n326 , n64 );
    or g522 ( n118 , n1148 , n1293 );
    xor g523 ( n1058 , n1060 , n171 );
    or g524 ( n1026 , n1213 , n1581 );
    or g525 ( n1055 , n1000 , n619 );
    and g526 ( n907 , n1259 , n593 );
    nor g527 ( n886 , n805 , n1320 );
    and g528 ( n1491 , n1644 , n752 );
    not g529 ( n518 , n480 );
    xnor g530 ( n993 , n50 , n1192 );
    or g531 ( n1150 , n149 , n1053 );
    nor g532 ( n10 , n555 , n927 );
    and g533 ( n756 , n155 , n1000 );
    not g534 ( n1300 , n1070 );
    not g535 ( n304 , n896 );
    xnor g536 ( n861 , n1636 , n1039 );
    and g537 ( n558 , n581 , n529 );
    not g538 ( n48 , n1639 );
    or g539 ( n808 , n920 , n1319 );
    and g540 ( n436 , n845 , n545 );
    and g541 ( n1137 , n41 , n844 );
    xnor g542 ( n619 , n508 , n379 );
    and g543 ( n1632 , n1643 , n761 );
    xnor g544 ( n1073 , n1307 , n480 );
    not g545 ( n1469 , n730 );
    not g546 ( n1615 , n162 );
    not g547 ( n720 , n1307 );
    not g548 ( n499 , n1187 );
    not g549 ( n21 , n691 );
    nor g550 ( n461 , n266 , n184 );
    xnor g551 ( n1340 , n745 , n1752 );
    not g552 ( n1696 , n1539 );
    not g553 ( n876 , n968 );
    and g554 ( n1148 , n1065 , n1598 );
    or g555 ( n578 , n1713 , n1443 );
    xnor g556 ( n1760 , n952 , n329 );
    or g557 ( n43 , n143 , n413 );
    nor g558 ( n1056 , n634 , n1357 );
    and g559 ( n111 , n1029 , n868 );
    or g560 ( n1404 , n300 , n28 );
    not g561 ( n1360 , n977 );
    nor g562 ( n15 , n1763 , n395 );
    not g563 ( n219 , n422 );
    nor g564 ( n835 , n410 , n1578 );
    and g565 ( n95 , n1149 , n1615 );
    and g566 ( n28 , n129 , n11 );
    xnor g567 ( n1736 , n1139 , n9 );
    and g568 ( n734 , n455 , n467 );
    or g569 ( n1124 , n815 , n281 );
    or g570 ( n1383 , n1388 , n907 );
    not g571 ( n1555 , n234 );
    or g572 ( n1014 , n1041 , n661 );
    or g573 ( n1110 , n337 , n30 );
    not g574 ( n564 , n542 );
    and g575 ( n383 , n687 , n83 );
    or g576 ( n404 , n926 , n1492 );
    not g577 ( n1744 , n1159 );
    or g578 ( n1297 , n652 , n78 );
    xnor g579 ( n792 , n153 , n1032 );
    and g580 ( n929 , n417 , n1019 );
    or g581 ( n1127 , n682 , n1371 );
    not g582 ( n406 , n1739 );
    xnor g583 ( n1113 , n849 , n898 );
    nor g584 ( n899 , n787 , n1280 );
    nor g585 ( n465 , n921 , n1549 );
    or g586 ( n1644 , n1750 , n582 );
    not g587 ( n1247 , n788 );
    not g588 ( n193 , n1418 );
    nor g589 ( n1640 , n562 , n993 );
    and g590 ( n770 , n35 , n1333 );
    not g591 ( n594 , n1003 );
    xnor g592 ( n1326 , n386 , n226 );
    or g593 ( n568 , n291 , n939 );
    not g594 ( n236 , n498 );
    xnor g595 ( n638 , n470 , n721 );
    not g596 ( n1180 , n1356 );
    nor g597 ( n1122 , n410 , n1560 );
    or g598 ( n806 , n1195 , n1581 );
    not g599 ( n437 , n1559 );
    and g600 ( n643 , n128 , n538 );
    or g601 ( n1177 , n1266 , n1612 );
    or g602 ( n985 , n926 , n562 );
    not g603 ( n1403 , n1658 );
    xnor g604 ( n1144 , n562 , n923 );
    or g605 ( n668 , n682 , n1000 );
    not g606 ( n1604 , n1045 );
    nor g607 ( n965 , n607 , n1678 );
    not g608 ( n358 , n801 );
    xnor g609 ( n1169 , n1034 , n637 );
    xnor g610 ( n966 , n353 , n498 );
    not g611 ( n369 , n171 );
    not g612 ( n1212 , n173 );
    or g613 ( n136 , n1381 , n89 );
    not g614 ( n716 , n818 );
    not g615 ( n964 , n1505 );
    or g616 ( n1431 , n1532 , n1163 );
    not g617 ( n1572 , n1610 );
    not g618 ( n1359 , n1409 );
    or g619 ( n571 , n1527 , n61 );
    not g620 ( n257 , n1033 );
    not g621 ( n732 , n1073 );
    not g622 ( n186 , n841 );
    xnor g623 ( n1021 , n353 , n695 );
    and g624 ( n301 , n1157 , n1190 );
    or g625 ( n1141 , n1640 , n451 );
    not g626 ( n1004 , n497 );
    xnor g627 ( n334 , n1082 , n37 );
    or g628 ( n29 , n1410 , n1612 );
    or g629 ( n1754 , n1123 , n249 );
    xnor g630 ( n290 , n1171 , n594 );
    or g631 ( n1290 , n1585 , n42 );
    or g632 ( n1444 , n379 , n709 );
    xnor g633 ( n216 , n894 , n1128 );
    or g634 ( n1132 , n556 , n1745 );
    not g635 ( n856 , n1655 );
    or g636 ( n954 , n757 , n348 );
    or g637 ( n1771 , n744 , n1031 );
    or g638 ( n1311 , n369 , n1167 );
    or g639 ( n1400 , n1266 , n407 );
    or g640 ( n844 , n1294 , n525 );
    or g641 ( n1107 , n1607 , n1536 );
    not g642 ( n565 , n435 );
    xnor g643 ( n979 , n1646 , n755 );
    not g644 ( n57 , n862 );
    not g645 ( n1203 , n714 );
    xnor g646 ( n1723 , n191 , n966 );
    not g647 ( n552 , n1591 );
    xnor g648 ( n75 , n528 , n1592 );
    and g649 ( n531 , n1674 , n420 );
    or g650 ( n988 , n1476 , n1491 );
    or g651 ( n1224 , n1263 , n1548 );
    and g652 ( n180 , n115 , n356 );
    or g653 ( n318 , n1146 , n1496 );
    xnor g654 ( n1409 , n1607 , n183 );
    xnor g655 ( n1629 , n383 , n1325 );
    not g656 ( n99 , n249 );
    not g657 ( n1266 , n1740 );
    or g658 ( n5 , n220 , n398 );
    and g659 ( n838 , n158 , n1406 );
    xnor g660 ( n1660 , n1391 , n793 );
    not g661 ( n1628 , n684 );
    or g662 ( n897 , n1758 , n1243 );
    or g663 ( n1693 , n166 , n1168 );
    or g664 ( n501 , n973 , n915 );
    and g665 ( n884 , n1597 , n1512 );
    not g666 ( n201 , n1274 );
    nor g667 ( n874 , n444 , n977 );
    or g668 ( n1638 , n697 , n1331 );
    or g669 ( n1088 , n1532 , n189 );
    nor g670 ( n357 , n1678 , n402 );
    nor g671 ( n513 , n693 , n1365 );
    and g672 ( n354 , n754 , n1557 );
    not g673 ( n1208 , n1104 );
    or g674 ( n1085 , n509 , n1013 );
    not g675 ( n127 , n17 );
    not g676 ( n1645 , n582 );
    and g677 ( n93 , n1744 , n1361 );
    nor g678 ( n556 , n555 , n788 );
    nor g679 ( n605 , n629 , n713 );
    not g680 ( n1513 , n26 );
    or g681 ( n958 , n310 , n1551 );
    or g682 ( n1233 , n1246 , n678 );
    or g683 ( n1406 , n1000 , n1131 );
    and g684 ( n280 , n1626 , n1164 );
    and g685 ( n603 , n257 , n1725 );
    or g686 ( n1571 , n105 , n881 );
    not g687 ( n1607 , n1145 );
    not g688 ( n1195 , n1070 );
    not g689 ( n576 , n633 );
    nor g690 ( n384 , n1196 , n1236 );
    and g691 ( n480 , n666 , n1749 );
    and g692 ( n1658 , n1237 , n1609 );
    not g693 ( n143 , n46 );
    or g694 ( n1545 , n650 , n134 );
    xnor g695 ( n242 , n104 , n1770 );
    and g696 ( n1745 , n1080 , n1286 );
    xnor g697 ( n238 , n1019 , n645 );
    nor g698 ( n864 , n1259 , n436 );
    and g699 ( n1450 , n956 , n1445 );
    xnor g700 ( n1521 , n879 , n679 );
    nor g701 ( n314 , n1341 , n1014 );
    and g702 ( n1691 , n607 , n266 );
    xnor g703 ( n1191 , n1664 , n58 );
    xnor g704 ( n1748 , n16 , n324 );
    or g705 ( n1439 , n885 , n539 );
    or g706 ( n288 , n742 , n1002 );
    not g707 ( n142 , n1221 );
    and g708 ( n79 , n870 , n1000 );
    or g709 ( n1692 , n359 , n636 );
    not g710 ( n1265 , n1213 );
    xnor g711 ( n1315 , n1727 , n1619 );
    or g712 ( n495 , n399 , n1205 );
    or g713 ( n2 , n614 , n364 );
    xnor g714 ( n1299 , n413 , n1320 );
    xnor g715 ( n677 , n1584 , n223 );
    xnor g716 ( n1283 , n1725 , n1494 );
    nor g717 ( n549 , n821 , n53 );
    or g718 ( n505 , n362 , n663 );
    nor g719 ( n918 , n1160 , n1532 );
    not g720 ( n543 , n1422 );
    not g721 ( n1167 , n266 );
    or g722 ( n162 , n1083 , n87 );
    or g723 ( n455 , n1225 , n1578 );
    not g724 ( n1742 , n692 );
    xnor g725 ( n905 , n1054 , n334 );
    not g726 ( n1387 , n628 );
    xnor g727 ( n405 , n1576 , n435 );
    nor g728 ( n850 , n1173 , n791 );
    or g729 ( n3 , n1597 , n1512 );
    not g730 ( n983 , n1288 );
    not g731 ( n364 , n580 );
    xnor g732 ( n488 , n166 , n347 );
    and g733 ( n184 , n1583 , n61 );
    and g734 ( n593 , n845 , n1421 );
    and g735 ( n647 , n962 , n1703 );
    or g736 ( n1231 , n1229 , n1563 );
    not g737 ( n289 , n414 );
    or g738 ( n1508 , n237 , n710 );
    or g739 ( n1206 , n562 , n713 );
    or g740 ( n385 , n1122 , n625 );
    or g741 ( n244 , n1670 , n1336 );
    xnor g742 ( n787 , n1732 , n839 );
    or g743 ( n1274 , n1513 , n1313 );
    not g744 ( n37 , n1164 );
    xnor g745 ( n1727 , n504 , n495 );
    not g746 ( n389 , n144 );
    not g747 ( n671 , n1022 );
    or g748 ( n1458 , n617 , n1719 );
    xnor g749 ( n658 , n1448 , n411 );
    or g750 ( n637 , n735 , n448 );
    and g751 ( n596 , n999 , n1517 );
    nor g752 ( n1309 , n703 , n604 );
    not g753 ( n1083 , n1731 );
    not g754 ( n1186 , n1111 );
    xnor g755 ( n1581 , n504 , n1228 );
    and g756 ( n763 , n1431 , n176 );
    xnor g757 ( n836 , n552 , n694 );
    not g758 ( n1250 , n504 );
    xnor g759 ( n423 , n1007 , n751 );
    xnor g760 ( n1142 , n1221 , n660 );
    not g761 ( n1017 , n1496 );
    or g762 ( n506 , n1123 , n1134 );
    xnor g763 ( n728 , n713 , n629 );
    and g764 ( n168 , n486 , n268 );
    not g765 ( n1443 , n977 );
    xnor g766 ( n712 , n1519 , n919 );
    nor g767 ( n624 , n1643 , n1707 );
    nor g768 ( n81 , n952 , n653 );
    and g769 ( n1278 , n1413 , n793 );
    not g770 ( n634 , n1109 );
    or g771 ( n774 , n577 , n1289 );
    and g772 ( n609 , n43 , n1772 );
    not g773 ( n1577 , n1172 );
    or g774 ( n25 , n962 , n160 );
    xnor g775 ( n1766 , n1208 , n1612 );
    xnor g776 ( n123 , n1745 , n785 );
    xnor g777 ( n419 , n816 , n968 );
    or g778 ( n206 , n820 , n402 );
    and g779 ( n187 , n205 , n225 );
    or g780 ( n1269 , n252 , n400 );
    or g781 ( n417 , n613 , n679 );
    or g782 ( n719 , n730 , n1186 );
    or g783 ( n85 , n1711 , n566 );
    or g784 ( n765 , n22 , n1477 );
    nor g785 ( n520 , n1371 , n716 );
    xnor g786 ( n698 , n1545 , n779 );
    not g787 ( n1232 , n544 );
    xnor g788 ( n491 , n1709 , n1643 );
    xnor g789 ( n1686 , n869 , n1681 );
    or g790 ( n1028 , n1636 , n1209 );
    not g791 ( n1134 , n729 );
    or g792 ( n8 , n1542 , n1773 );
    not g793 ( n1683 , n617 );
    not g794 ( n224 , n1623 );
    nor g795 ( n1294 , n1512 , n271 );
    or g796 ( n411 , n1603 , n1291 );
    or g797 ( n821 , n1673 , n843 );
    xnor g798 ( n1498 , n1289 , n1395 );
    nor g799 ( n1006 , n1264 , n524 );
    not g800 ( n537 , n1433 );
    nor g801 ( n134 , n1066 , n1614 );
    or g802 ( n978 , n291 , n1366 );
    not g803 ( n1045 , n900 );
    or g804 ( n467 , n168 , n311 );
    xnor g805 ( n1330 , n1396 , n686 );
    or g806 ( n956 , n1751 , n1226 );
    not g807 ( n666 , n1575 );
    nor g808 ( n310 , n1263 , n483 );
    xnor g809 ( n489 , n173 , n1501 );
    xnor g810 ( n58 , n362 , n374 );
    xnor g811 ( n919 , n1473 , n791 );
    nor g812 ( n1514 , n257 , n261 );
    nor g813 ( n355 , n926 , n211 );
    not g814 ( n569 , n20 );
    not g815 ( n1506 , n50 );
    or g816 ( n340 , n1151 , n671 );
    xnor g817 ( n67 , n1653 , n214 );
    and g818 ( n1549 , n531 , n1446 );
    not g819 ( n365 , n1490 );
    or g820 ( n877 , n730 , n373 );
    and g821 ( n333 , n212 , n1587 );
    or g822 ( n633 , n1702 , n445 );
    xnor g823 ( n755 , n1300 , n298 );
    xnor g824 ( n243 , n265 , n952 );
    not g825 ( n937 , n1434 );
    and g826 ( n997 , n1520 , n1016 );
    xnor g827 ( n1202 , n647 , n646 );
    xnor g828 ( n476 , n1071 , n1069 );
    not g829 ( n674 , n265 );
    xnor g830 ( n1235 , n1364 , n719 );
    xnor g831 ( n779 , n1371 , n682 );
    not g832 ( n297 , n600 );
    xnor g833 ( n172 , n1230 , n602 );
    and g834 ( n1625 , n1464 , n1200 );
    or g835 ( n793 , n567 , n1074 );
    nor g836 ( n1178 , n353 , n1351 );
    xnor g837 ( n950 , n1612 , n722 );
    or g838 ( n1252 , n1607 , n893 );
    nor g839 ( n1196 , n164 , n682 );
    xnor g840 ( n547 , n691 , n1718 );
    xnor g841 ( n372 , n83 , n1189 );
    not g842 ( n1687 , n1450 );
    or g843 ( n1569 , n740 , n1389 );
    not g844 ( n799 , n656 );
    or g845 ( n1470 , n77 , n1421 );
    xnor g846 ( n156 , n1602 , n342 );
    nor g847 ( n279 , n464 , n1007 );
    not g848 ( n137 , n254 );
    or g849 ( n776 , n899 , n550 );
    not g850 ( n1656 , n539 );
    and g851 ( n430 , n869 , n470 );
    or g852 ( n566 , n266 , n1471 );
    and g853 ( n606 , n86 , n592 );
    or g854 ( n341 , n226 , n386 );
    not g855 ( n1248 , n346 );
    and g856 ( n986 , n1223 , n553 );
    xnor g857 ( n270 , n1364 , n877 );
    or g858 ( n502 , n1114 , n705 );
    xnor g859 ( n1325 , n1253 , n1031 );
    not g860 ( n483 , n1548 );
    and g861 ( n1022 , n1687 , n1424 );
    not g862 ( n893 , n931 );
    xnor g863 ( n1405 , n1456 , n783 );
    not g864 ( n775 , n996 );
    not g865 ( n805 , n163 );
    or g866 ( n1772 , n443 , n880 );
    and g867 ( n736 , n742 , n1503 );
    nor g868 ( n399 , n1275 , n18 );
    xnor g869 ( n1194 , n1118 , n1087 );
    not g870 ( n24 , n1405 );
    or g871 ( n1386 , n1390 , n463 );
    not g872 ( n1357 , n281 );
    xnor g873 ( n74 , n983 , n1630 );
    or g874 ( n631 , n662 , n1625 );
    and g875 ( n1636 , n767 , n345 );
    not g876 ( n377 , n1678 );
    nor g877 ( n120 , n241 , n100 );
    or g878 ( n1276 , n1350 , n1303 );
    xnor g879 ( n1185 , n331 , n606 );
    xnor g880 ( n626 , n936 , n1530 );
    or g881 ( n718 , n1426 , n96 );
    nor g882 ( n853 , n1174 , n37 );
    xnor g883 ( n429 , n873 , n493 );
    xnor g884 ( n1733 , n490 , n1335 );
    nor g885 ( n746 , n132 , n383 );
    xnor g886 ( n1553 , n1575 , n1490 );
    xnor g887 ( n1677 , n570 , n419 );
    and g888 ( n1214 , n1537 , n896 );
    xnor g889 ( n1601 , n1614 , n521 );
    xnor g890 ( n721 , n441 , n1539 );
    not g891 ( n1706 , n940 );
    nor g892 ( n199 , n164 , n968 );
    not g893 ( n164 , n402 );
    and g894 ( n550 , n29 , n546 );
    xnor g895 ( n969 , n1623 , n799 );
    or g896 ( n267 , n349 , n714 );
    and g897 ( n396 , n449 , n32 );
    not g898 ( n1354 , n400 );
    nor g899 ( n89 , n583 , n1092 );
    xnor g900 ( n1731 , n326 , n1227 );
    xnor g901 ( n1237 , n633 , n1145 );
    xnor g902 ( n181 , n960 , n1541 );
    xnor g903 ( n828 , n562 , n1221 );
    and g904 ( n1111 , n581 , n804 );
    and g905 ( n507 , n766 , n1559 );
    xnor g906 ( n645 , n679 , n613 );
    xnor g907 ( n790 , n525 , n1304 );
    or g908 ( n1345 , n1301 , n609 );
    not g909 ( n441 , n1427 );
    and g910 ( n650 , n1435 , n1174 );
    nor g911 ( n154 , n213 , n1360 );
    xnor g912 ( n1570 , n1626 , n37 );
    or g913 ( n1454 , n1254 , n903 );
    or g914 ( n1561 , n359 , n977 );
    not g915 ( n343 , n1222 );
    xnor g916 ( n486 , n519 , n649 );
    xnor g917 ( n694 , n1229 , n1031 );
    xnor g918 ( n1460 , n261 , n670 );
    xor g919 ( n1103 , n715 , n1565 );
    or g920 ( n933 , n1295 , n169 );
    not g921 ( n1270 , n228 );
    and g922 ( n1567 , n1181 , n1436 );
    xnor g923 ( n1012 , n1599 , n575 );
    not g924 ( n1192 , n301 );
    and g925 ( n970 , n834 , n481 );
    and g926 ( n282 , n1489 , n167 );
    and g927 ( n313 , n1026 , n988 );
    and g928 ( n533 , n1734 , n1639 );
    not g929 ( n1310 , n35 );
    or g930 ( n1618 , n918 , n1241 );
    or g931 ( n1541 , n718 , n698 );
    or g932 ( n1060 , n1768 , n871 );
    or g933 ( n221 , n471 , n152 );
    or g934 ( n1735 , n101 , n1167 );
    not g935 ( n1209 , n1002 );
    or g936 ( n1162 , n540 , n804 );
    not g937 ( n581 , n1118 );
    or g938 ( n1429 , n1123 , n1153 );
    nor g939 ( n207 , n1480 , n104 );
    or g940 ( n1548 , n379 , n571 );
    or g941 ( n1044 , n413 , n1405 );
    not g942 ( n1655 , n1401 );
    and g943 ( n681 , n1747 , n1455 );
    or g944 ( n245 , n291 , n1247 );
    xnor g945 ( n1654 , n1477 , n319 );
    and g946 ( n656 , n1238 , n872 );
    xnor g947 ( n1067 , n502 , n1106 );
    or g948 ( n119 , n737 , n1742 );
    xnor g949 ( n521 , n1174 , n1435 );
    not g950 ( n130 , n88 );
    or g951 ( n688 , n1253 , n1 );
    nor g952 ( n1710 , n47 , n1207 );
    nor g953 ( n875 , n1643 , n424 );
    and g954 ( n1288 , n1756 , n840 );
    not g955 ( n1016 , n1244 );
    xnor g956 ( n344 , n1643 , n469 );
    or g957 ( n1154 , n1632 , n984 );
    xnor g958 ( n630 , n1300 , n967 );
    and g959 ( n1380 , n1059 , n818 );
    and g960 ( n1500 , n1381 , n1697 );
    or g961 ( n225 , n1669 , n1579 );
    nor g962 ( n478 , n562 , n1664 );
    or g963 ( n16 , n913 , n461 );
    xnor g964 ( n117 , n490 , n1585 );
    and g965 ( n1519 , n1003 , n1171 );
    and g966 ( n1651 , n1027 , n1482 );
    or g967 ( n1008 , n161 , n187 );
    or g968 ( n772 , n1381 , n743 );
    or g969 ( n1157 , n838 , n1187 );
    or g970 ( n589 , n1178 , n320 );
    nor g971 ( n1066 , n1435 , n1174 );
    or g972 ( n1703 , n1145 , n275 );
    nor g973 ( n1102 , n1743 , n197 );
    xnor g974 ( n1348 , n128 , n538 );
    and g975 ( n1379 , n815 , n281 );
    nor g976 ( n1761 , n170 , n1762 );
    nor g977 ( n1377 , n69 , n98 );
    or g978 ( n356 , n479 , n375 );
    xnor g979 ( n1516 , n555 , n1363 );
    and g980 ( n1484 , n1341 , n1014 );
    not g981 ( n1104 , n1740 );
    and g982 ( n1187 , n656 , n224 );
    or g983 ( n723 , n820 , n1402 );
    and g984 ( n620 , n1561 , n1569 );
    or g985 ( n1218 , n1684 , n39 );
    or g986 ( n957 , n1160 , n1167 );
    nor g987 ( n450 , n369 , n402 );
    or g988 ( n62 , n1390 , n582 );
    and g989 ( n182 , n1497 , n1061 );
    nor g990 ( n107 , n90 , n513 );
    or g991 ( n1048 , n928 , n122 );
    or g992 ( n1559 , n909 , n107 );
    or g993 ( n151 , n442 , n1550 );
    xnor g994 ( n1305 , n35 , n907 );
    not g995 ( n796 , n757 );
    nor g996 ( n601 , n1130 , n1220 );
    and g997 ( n852 , n177 , n571 );
    xnor g998 ( n284 , n318 , n1159 );
    and g999 ( n1438 , n1461 , n1000 );
    or g1000 ( n1397 , n666 , n1193 );
    and g1001 ( n741 , n543 , n159 );
    xnor g1002 ( n1260 , n76 , n430 );
    or g1003 ( n152 , n428 , n258 );
    not g1004 ( n967 , n72 );
    or g1005 ( n1452 , n291 , n735 );
    not g1006 ( n519 , n1182 );
    and g1007 ( n504 , n1524 , n204 );
    not g1008 ( n97 , n1151 );
    nor g1009 ( n6 , n257 , n1382 );
    or g1010 ( n1337 , n1329 , n490 );
    or g1011 ( n833 , n1229 , n1693 );
    or g1012 ( n1554 , n359 , n802 );
    or g1013 ( n1433 , n1509 , n287 );
    and g1014 ( n1143 , n285 , n278 );
    xnor g1015 ( n1061 , n1418 , n1010 );
    or g1016 ( n360 , n410 , n400 );
    or g1017 ( n211 , n379 , n88 );
    xnor g1018 ( n1675 , n228 , n572 );
    xnor g1019 ( n753 , n16 , n114 );
    xnor g1020 ( n1415 , n596 , n1516 );
    not g1021 ( n447 , n889 );
    and g1022 ( n1671 , n1452 , n1378 );
    not g1023 ( n166 , n438 );
    not g1024 ( n608 , n91 );
    or g1025 ( n975 , n1266 , n602 );
    and g1026 ( n54 , n1631 , n668 );
    or g1027 ( n1002 , n16 , n1462 );
    not g1028 ( n804 , n1087 );
    and g1029 ( n23 , n422 , n1618 );
    xnor g1030 ( n1507 , n1319 , n1736 );
    or g1031 ( n999 , n359 , n236 );
    xnor g1032 ( n832 , n333 , n1668 );
    or g1033 ( n685 , n1380 , n425 );
    xnor g1034 ( n991 , n933 , n1098 );
    not g1035 ( n1442 , n1109 );
    and g1036 ( n1226 , n735 , n977 );
    or g1037 ( n1650 , n1379 , n651 );
    not g1038 ( n868 , n340 );
    and g1039 ( n1681 , n1206 , n385 );
    not g1040 ( n1109 , n612 );
    or g1041 ( n86 , n965 , n946 );
    or g1042 ( n962 , n1607 , n408 );
    xnor g1043 ( n72 , n1022 , n97 );
    xnor g1044 ( n239 , n952 , n729 );
    xnor g1045 ( n803 , n1448 , n555 );
    xnor g1046 ( n215 , n1371 , n1555 );
    or g1047 ( n538 , n1602 , n1297 );
    not g1048 ( n1382 , n1563 );
    xnor g1049 ( n1168 , n275 , n801 );
    xnor g1050 ( n1585 , n90 , n951 );
    or g1051 ( n1489 , n157 , n674 );
    not g1052 ( n1339 , n195 );
    or g1053 ( n632 , n1123 , n289 );
    xnor g1054 ( n1497 , n320 , n248 );
    not g1055 ( n185 , n1370 );
    not g1056 ( n373 , n558 );
    xnor g1057 ( n1139 , n375 , n1023 );
    xnor g1058 ( n1543 , n1468 , n537 );
    or g1059 ( n1591 , n166 , n849 );
    not g1060 ( n1536 , n183 );
    not g1061 ( n1534 , n1228 );
    nor g1062 ( n895 , n555 , n1363 );
    or g1063 ( n1728 , n800 , n323 );
    or g1064 ( n859 , n1195 , n298 );
    or g1065 ( n1052 , n266 , n784 );
    and g1066 ( n1095 , n720 , n178 );
    or g1067 ( n457 , n514 , n529 );
    or g1068 ( n1515 , n562 , n386 );
    xnor g1069 ( n1505 , n970 , n368 );
    nor g1070 ( n984 , n1682 , n180 );
    not g1071 ( n679 , n1553 );
    or g1072 ( n1605 , n854 , n929 );
    xnor g1073 ( n1373 , n1750 , n1645 );
    not g1074 ( n255 , n847 );
    or g1075 ( n1436 , n1362 , n831 );
    or g1076 ( n1240 , n198 , n1308 );
    xnor g1077 ( n1538 , n1266 , n39 );
    or g1078 ( n1575 , n925 , n717 );
    xnor g1079 ( n1653 , n389 , n608 );
    or g1080 ( n1518 , n82 , n1334 );
    xnor g1081 ( n912 , n1118 , n119 );
    or g1082 ( n657 , n1266 , n861 );
    not g1083 ( n1680 , n1227 );
    xnor g1084 ( n386 , n652 , n346 );
    or g1085 ( n294 , n814 , n1562 );
    xnor g1086 ( n683 , n1150 , n1081 );
    and g1087 ( n1419 , n1218 , n1150 );
    and g1088 ( n544 , n820 , n1402 );
    xnor g1089 ( n1573 , n1643 , n424 );
    or g1090 ( n210 , n150 , n1441 );
    or g1091 ( n1635 , n1649 , n250 );
    or g1092 ( n265 , n492 , n976 );
    xnor g1093 ( n1672 , n396 , n1434 );
    or g1094 ( n1007 , n1047 , n850 );
    not g1095 ( n1256 , n156 );
    and g1096 ( n706 , n985 , n1233 );
    xnor g1097 ( n771 , n764 , n170 );
    or g1098 ( n990 , n1256 , n1487 );
    nor g1099 ( n1648 , n926 , n1548 );
    not g1100 ( n1423 , n870 );
    not g1101 ( n1599 , n1011 );
    not g1102 ( n163 , n307 );
    and g1103 ( n1198 , n325 , n380 );
    not g1104 ( n865 , n306 );
    or g1105 ( n1416 , n1282 , n234 );
    or g1106 ( n872 , n1000 , n388 );
    not g1107 ( n1713 , n444 );
    xnor g1108 ( n1176 , n555 , n927 );
    xnor g1109 ( n1131 , n293 , n1422 );
    not g1110 ( n816 , n515 );
    nor g1111 ( n615 , n155 , n402 );
    nor g1112 ( n1344 , n353 , n747 );
    or g1113 ( n87 , n284 , n2 );
    nor g1114 ( n1689 , n379 , n1217 );
    and g1115 ( n977 , n109 , n192 );
    not g1116 ( n410 , n889 );
    or g1117 ( n1447 , n1285 , n371 );
    buf g1118 ( n1217 , n1712 );
    or g1119 ( n940 , n1597 , n682 );
    not g1120 ( n453 , n1240 );
    not g1121 ( n1329 , n66 );
    nor g1122 ( n1170 , n1208 , n39 );
    or g1123 ( n335 , n369 , n1060 );
    xnor g1124 ( n1408 , n1651 , n491 );
    xnor g1125 ( n690 , n1706 , n46 );
    nor g1126 ( n1704 , n1466 , n745 );
    not g1127 ( n760 , n1549 );
    xnor g1128 ( n1101 , n26 , n607 );
    xnor g1129 ( n139 , n562 , n1312 );
    nor g1130 ( n1246 , n1263 , n447 );
    and g1131 ( n1287 , n1673 , n1079 );
    not g1132 ( n1411 , n49 );
    and g1133 ( n232 , n40 , n75 );
    not g1134 ( n1171 , n626 );
    and g1135 ( n660 , n663 , n1753 );
    not g1136 ( n1468 , n528 );
    or g1137 ( n955 , n1123 , n674 );
    or g1138 ( n1424 , n1608 , n496 );
    xnor g1139 ( n401 , n190 , n950 );
    or g1140 ( n992 , n280 , n817 );
    not g1141 ( n560 , n747 );
    or g1142 ( n691 , n1621 , n1368 );
    xnor g1143 ( n378 , n1662 , n328 );
    not g1144 ( n38 , n1204 );
    and g1145 ( n892 , n1413 , n1755 );
    and g1146 ( n1009 , n143 , n1285 );
    xnor g1147 ( n471 , n1636 , n246 );
    or g1148 ( n1587 , n1377 , n282 );
    nor g1149 ( n418 , n952 , n329 );
    xnor g1150 ( n286 , n1672 , n1217 );
    xnor g1151 ( n914 , n1428 , n239 );
    xnor g1152 ( n848 , n353 , n747 );
    xnor g1153 ( n1057 , n45 , n1573 );
    or g1154 ( n1767 , n1056 , n639 );
    nor g1155 ( n1529 , n1643 , n469 );
    and g1156 ( n831 , n1465 , n685 );
    or g1157 ( n1020 , n207 , n847 );
    nor g1158 ( n784 , n177 , n571 );
    not g1159 ( n327 , n655 );
    not g1160 ( n782 , n1616 );
    xnor g1161 ( n426 , n1243 , n1701 );
    or g1162 ( n251 , n6 , n1579 );
    xnor g1163 ( n930 , n952 , n1296 );
    not g1164 ( n114 , n466 );
    or g1165 ( n446 , n1219 , n1553 );
    xnor g1166 ( n559 , n434 , n405 );
    xnor g1167 ( n1480 , n916 , n906 );
    not g1168 ( n644 , n1198 );
    nor g1169 ( n1758 , n1174 , n9 );
    or g1170 ( n256 , n413 , n753 );
    xnor g1171 ( n179 , n1594 , n1430 );
    or g1172 ( n459 , n884 , n421 );
    not g1173 ( n1328 , n1332 );
    or g1174 ( n115 , n291 , n1577 );
    and g1175 ( n579 , n1195 , n298 );
    and g1176 ( n1074 , n1515 , n1522 );
    xnor g1177 ( n1395 , n1415 , n351 );
    xnor g1178 ( n942 , n152 , n1119 );
    xnor g1179 ( n1175 , n221 , n865 );
    not g1180 ( n296 , n1313 );
    or g1181 ( n1531 , n1381 , n811 );
    not g1182 ( n1 , n383 );
    or g1183 ( n1394 , n362 , n142 );
    not g1184 ( n1336 , n1528 );
    not g1185 ( n1136 , n972 );
    nor g1186 ( n1205 , n590 , n1651 );
    nor g1187 ( n1350 , n1512 , n967 );
    not g1188 ( n1532 , n1000 );
    not g1189 ( n463 , n1169 );
    xnor g1190 ( n1737 , n76 , n53 );
    and g1191 ( n320 , n506 , n1036 );
    nor g1192 ( n1590 , n1422 , n230 );
    xnor g1193 ( n1282 , n370 , n344 );
    nor g1194 ( n262 , n353 , n695 );
    or g1195 ( n1027 , n291 , n523 );
    buf g1196 ( n1712 , n1314 );
    or g1197 ( n1434 , n465 , n224 );
    xnor g1198 ( n981 , n1497 , n1335 );
    not g1199 ( n567 , n1165 );
    or g1200 ( n1163 , n866 , n201 );
    or g1201 ( n598 , n1392 , n1273 );
    xnor g1202 ( n468 , n1059 , n716 );
    or g1203 ( n910 , n235 , n143 );
    xnor g1204 ( n699 , n1188 , n1144 );
    or g1205 ( n1117 , n1720 , n635 );
    xnor g1206 ( n1600 , n943 , n1451 );
    or g1207 ( n92 , n1602 , n1716 );
    nor g1208 ( n1682 , n1643 , n761 );
    xnor g1209 ( n218 , n187 , n381 );
    not g1210 ( n350 , n1681 );
    not g1211 ( n440 , n1764 );
    and g1212 ( n1041 , n155 , n1381 );
    and g1213 ( n1708 , n1088 , n393 );
    or g1214 ( n1652 , n914 , n798 );
    and g1215 ( n841 , n606 , n1647 );
    xnor g1216 ( n1698 , n1582 , n967 );
    xnor g1217 ( n1630 , n1555 , n1634 );
    xnor g1218 ( n1128 , n40 , n271 );
    nor g1219 ( n794 , n1527 , n1009 );
    nor g1220 ( n309 , n607 , n402 );
    and g1221 ( n105 , n952 , n653 );
    or g1222 ( n233 , n20 , n1458 );
    xnor g1223 ( n403 , n584 , n1560 );
    or g1224 ( n1448 , n1540 , n938 );
    and g1225 ( n972 , n1028 , n288 );
    and g1226 ( n909 , n693 , n1365 );
    not g1227 ( n1229 , n515 );
    or g1228 ( n1623 , n778 , n760 );
    or g1229 ( n526 , n1586 , n1356 );
    not g1230 ( n879 , n1712 );
    not g1231 ( n1189 , n687 );
    xnor g1232 ( n517 , n1550 , n1521 );
    xnor g1233 ( n686 , n1672 , n1065 );
    xnor g1234 ( n1495 , n595 , n981 );
    xnor g1235 ( n381 , n1723 , n964 );
    and g1236 ( n1356 , n762 , n776 );
    or g1237 ( n752 , n702 , n1239 );
    xnor g1238 ( n1718 , n490 , n66 );
    or g1239 ( n1428 , n1607 , n1628 );
    and g1240 ( n1105 , n1751 , n1226 );
    xnor g1241 ( n317 , n313 , n771 );
    nor g1242 ( n427 , n1529 , n370 );
    not g1243 ( n494 , n1095 );
    or g1244 ( n503 , n413 , n435 );
    xnor g1245 ( n281 , n282 , n1267 );
    not g1246 ( n778 , n921 );
    or g1247 ( n397 , n358 , n408 );
    or g1248 ( n272 , n297 , n408 );
    nor g1249 ( n1241 , n876 , n1000 );
    or g1250 ( n701 , n116 , n1288 );
    and g1251 ( n191 , n632 , n945 );
    or g1252 ( n109 , n1423 , n1167 );
    not g1253 ( n636 , n1351 );
    and g1254 ( n1485 , n961 , n1387 );
    xnor g1255 ( n31 , n1643 , n36 );
    or g1256 ( n34 , n1219 , n1284 );
    xnor g1257 ( n614 , n911 , n1017 );
    not g1258 ( n302 , n986 );
    not g1259 ( n1487 , n95 );
    and g1260 ( n591 , n1183 , n1457 );
    nor g1261 ( n661 , n1417 , n830 );
    not g1262 ( n766 , n1120 );
    xnor g1263 ( n231 , n467 , n1475 );
    and g1264 ( n1093 , n1355 , n71 );
    or g1265 ( n1051 , n756 , n1449 );
    and g1266 ( n934 , n38 , n561 );
    not g1267 ( n1275 , n1643 );
    xnor g1268 ( n259 , n99 , n952 );
    and g1269 ( n150 , n1643 , n424 );
    not g1270 ( n553 , n458 );
    or g1271 ( n923 , n120 , n669 );
    or g1272 ( n1510 , n1607 , n1637 );
    or g1273 ( n908 , n306 , n221 );
    or g1274 ( n1738 , n1689 , n542 );
    or g1275 ( n1755 , n567 , n707 );
    not g1276 ( n348 , n507 );
    and g1277 ( n1562 , n1127 , n1545 );
    and g1278 ( n421 , n3 , n294 );
    or g1279 ( n1631 , n1532 , n1678 );
    and g1280 ( n1303 , n512 , n1412 );
    and g1281 ( n707 , n341 , n526 );
    nor g1282 ( n881 , n1437 , n81 );
    and g1283 ( n1402 , n1513 , n530 );
    xnor g1284 ( n439 , n628 , n961 );
    not g1285 ( n1108 , n1724 );
    and g1286 ( n1396 , n664 , n1020 );
    not g1287 ( n789 , n1743 );
    xnor g1288 ( n960 , n294 , n941 );
    xnor g1289 ( n904 , n439 , n753 );
    xnor g1290 ( n751 , n1585 , n1542 );
    not g1291 ( n175 , n69 );
    nor g1292 ( n621 , n450 , n750 );
    not g1293 ( n791 , n1398 );
    nor g1294 ( n1152 , n164 , n1597 );
    and g1295 ( n1307 , n1311 , n958 );
    or g1296 ( n1158 , n164 , n768 );
    or g1297 ( n141 , n330 , n764 );
    not g1298 ( n1446 , n412 );
    not g1299 ( n1624 , n159 );
    not g1300 ( n713 , n1560 );
    and g1301 ( n887 , n1527 , n1009 );
    not g1302 ( n1335 , n1061 );
    or g1303 ( n1679 , n876 , n266 );
    or g1304 ( n725 , n997 , n1719 );
    nor g1305 ( n982 , n667 , n1000 );
    xnor g1306 ( n1244 , n1389 , n812 );
    xnor g1307 ( n298 , n1185 , n954 );
    or g1308 ( n128 , n148 , n1500 );
    not g1309 ( n1123 , n952 );
    or g1310 ( n1200 , n1358 , n943 );
    xnor g1311 ( n610 , n1354 , n165 );
    or g1312 ( n1238 , n1532 , n1058 );
    and g1313 ( n1159 , n1596 , n146 );
    and g1314 ( n1227 , n1744 , n394 );
    and g1315 ( n651 , n688 , n1097 );
    xnor g1316 ( n867 , n392 , n1538 );
    and g1317 ( n161 , n1723 , n1505 );
    or g1318 ( n994 , n603 , n59 );
    xnor g1319 ( n823 , n651 , n1730 );
    not g1320 ( n1421 , n877 );
    nor g1321 ( n822 , n952 , n414 );
    nor g1322 ( n769 , n472 , n197 );
    nor g1323 ( n739 , n200 , n73 );
    nor g1324 ( n240 , n555 , n1448 );
    or g1325 ( n331 , n641 , n1420 );
    not g1326 ( n101 , n557 );
    xnor g1327 ( n1221 , n70 , n51 );
    not g1328 ( n1086 , n609 );
    nor g1329 ( n878 , n562 , n1221 );
    or g1330 ( n1522 , n321 , n1546 );
    not g1331 ( n1390 , n1045 );
    and g1332 ( n1207 , n245 , n1132 );
    nor g1333 ( n1301 , n1527 , n1208 );
    nor g1334 ( n697 , n634 , n964 );
    not g1335 ( n4 , n602 );
    and g1336 ( n388 , n404 , n696 );
    and g1337 ( n252 , n277 , n1376 );
    nor g1338 ( n1441 , n875 , n45 );
    xnor g1339 ( n1049 , n362 , n400 );
    not g1340 ( n508 , n709 );
    xnor g1341 ( n435 , n1748 , n340 );
    nor g1342 ( n299 , n821 , n430 );
    xnor g1343 ( n1494 , n257 , n1398 );
    xnor g1344 ( n91 , n441 , n264 );
    xnor g1345 ( n1633 , n1467 , n274 );
    xnor g1346 ( n1253 , n1510 , n930 );
    or g1347 ( n1096 , n1514 , n138 );
    xnor g1348 ( n1740 , n304 , n1537 );
    not g1349 ( n178 , n1397 );
    or g1350 ( n1375 , n54 , n1268 );
    and g1351 ( n1273 , n642 , n897 );
    nor g1352 ( n1649 , n1665 , n1667 );
    or g1353 ( n1039 , n366 , n466 );
    nor g1354 ( n59 , n1589 , n791 );
    and g1355 ( n896 , n433 , n1342 );
    or g1356 ( n936 , n1438 , n982 );
    nor g1357 ( n623 , n314 , n333 );
    not g1358 ( n1298 , n210 );
    or g1359 ( n1306 , n1381 , n1035 );
    xnor g1360 ( n1701 , n825 , n9 );
    xnor g1361 ( n588 , n625 , n403 );
    or g1362 ( n1188 , n878 , n1001 );
    and g1363 ( n625 , n446 , n151 );
    or g1364 ( n167 , n454 , n1759 );
    xnor g1365 ( n328 , n1734 , n48 );
    or g1366 ( n1619 , n1408 , n527 );
    xnor g1367 ( n276 , n1210 , n689 );
    xnor g1368 ( n1166 , n562 , n1263 );
    or g1369 ( n332 , n1245 , n113 );
    and g1370 ( n574 , n910 , n88 );
    nor g1371 ( n140 , n1601 , n1667 );
    or g1372 ( n1557 , n484 , n1198 );
    and g1373 ( n920 , n1139 , n832 );
    nor g1374 ( n1125 , n952 , n729 );
    not g1375 ( n1493 , n1455 );
    xnor g1376 ( n1746 , n635 , n376 );
    xnor g1377 ( n812 , n1443 , n353 );
    xnor g1378 ( n842 , n1770 , n1527 );
    nor g1379 ( n253 , n439 , n1320 );
    or g1380 ( n159 , n1263 , n211 );
    and g1381 ( n703 , n879 , n1672 );
    not g1382 ( n959 , n1214 );
    and g1383 ( n1343 , n876 , n570 );
    xnor g1384 ( n1338 , n1303 , n630 );
    and g1385 ( n1751 , n1478 , n963 );
    and g1386 ( n1490 , n742 , n1726 );
    or g1387 ( n1464 , n1082 , n658 );
    and g1388 ( n527 , n680 , n1739 );
    or g1389 ( n1076 , n1705 , n1318 );
    xnor g1390 ( n1025 , n374 , n1272 );
    or g1391 ( n285 , n1339 , n435 );
    not g1392 ( n783 , n973 );
    not g1393 ( n509 , n612 );
    not g1394 ( n1285 , n1597 );
    xnor g1395 ( n1481 , n1353 , n898 );
    nor g1396 ( n1264 , n164 , n46 );
    not g1397 ( n1071 , n1168 );
    not g1398 ( n1374 , n98 );
    or g1399 ( n1271 , n1078 , n873 );
    or g1400 ( n1190 , n339 , n499 );
    not g1401 ( n315 , n652 );
    xnor g1402 ( n1626 , n1318 , n409 );
    not g1403 ( n261 , n1693 );
    and g1404 ( n652 , n84 , n672 );
    nor g1405 ( n475 , n374 , n1179 );
    and g1406 ( n324 , n1468 , n1105 );
    or g1407 ( n1610 , n1258 , n427 );
    xnor g1408 ( n622 , n1643 , n761 );
    xnor g1409 ( n464 , n1571 , n786 );
    not g1410 ( n490 , n612 );
    not g1411 ( n197 , n249 );
    nor g1412 ( n1043 , n805 , n24 );
    or g1413 ( n532 , n1292 , n545 );
    and g1414 ( n337 , n1266 , n1612 );
    not g1415 ( n1466 , n914 );
    xnor g1416 ( n1399 , n1382 , n726 );
    xnor g1417 ( n138 , n397 , n1077 );
    and g1418 ( n1603 , n213 , n1360 );
    not g1419 ( n562 , n856 );
    and g1420 ( n1075 , n859 , n932 );
    and g1421 ( n894 , n485 , n1518 );
    nor g1422 ( n837 , n1230 , n4 );
    or g1423 ( n1228 , n18 , n217 );
    xnor g1424 ( n1568 , n1610 , n49 );
    not g1425 ( n880 , n459 );
    not g1426 ( n1462 , n324 );
    xnor g1427 ( n1078 , n441 , n1095 );
    xnor g1428 ( n1267 , n98 , n69 );
    and g1429 ( n1258 , n1643 , n469 );
    not g1430 ( n939 , n1140 );
    nor g1431 ( n1705 , n555 , n1140 );
    xnor g1432 ( n19 , n196 , n1262 );
    or g1433 ( n275 , n147 , n1091 );
    xnor g1434 ( n1033 , n1252 , n1760 );
    or g1435 ( n1236 , n1381 , n357 );
    nor g1436 ( n1504 , n1576 , n565 );
    not g1437 ( n1646 , n354 );
    xnor g1438 ( n1314 , n959 , n675 );
    xnor g1439 ( n737 , n459 , n890 );
    not g1440 ( n795 , n1581 );
    or g1441 ( n380 , n1384 , n13 );
    xnor g1442 ( n1535 , n817 , n1570 );
    xnor g1443 ( n1668 , n1014 , n1341 );
    and g1444 ( n1042 , n1211 , n1050 );
    nor g1445 ( n492 , n1160 , n1316 );
    or g1446 ( n1080 , n359 , n560 );
    xnor g1447 ( n941 , n1512 , n1597 );
    not g1448 ( n1721 , n680 );
    not g1449 ( n27 , n1485 );
    xnor g1450 ( n722 , n487 , n1757 );
    or g1451 ( n133 , n1427 , n1696 );
    or g1452 ( n1474 , n1484 , n623 );
    or g1453 ( n1024 , n235 , n782 );
    not g1454 ( n94 , n781 );
    and g1455 ( n1662 , n8 , n1279 );
    and g1456 ( n1526 , n379 , n130 );
    not g1457 ( n1371 , n900 );
    xnor g1458 ( n813 , n1334 , n1302 );
    or g1459 ( n1574 , n52 , n63 );
    and g1460 ( n577 , n1415 , n658 );
    nor g1461 ( n116 , n1634 , n1555 );
    xnor g1462 ( n1059 , n1147 , n1046 );
    nor g1463 ( n855 , n1643 , n1034 );
    or g1464 ( n592 , n1000 , n1094 );
    not g1465 ( n1670 , n1287 );
    xnor g1466 ( n135 , n425 , n468 );
    not g1467 ( n359 , n353 );
    and g1468 ( n1666 , n1643 , n36 );
    or g1469 ( n1197 , n164 , n1526 );
    and g1470 ( n392 , n256 , n1133 );
    or g1471 ( n1215 , n5 , n15 );
    or g1472 ( n60 , n1704 , n138 );
    xnor g1473 ( n1277 , n908 , n1249 );
    xnor g1474 ( n1164 , n1216 , n677 );
    and g1475 ( n1413 , n128 , n92 );
    not g1476 ( n330 , n170 );
    not g1477 ( n545 , n719 );
    not g1478 ( n1219 , n1712 );
    nor g1479 ( n885 , n781 , n24 );
    nor g1480 ( n563 , n164 , n66 );
    not g1481 ( n220 , n1530 );
    xnor g1482 ( n195 , n810 , n391 );
    and g1483 ( n1179 , n584 , n1664 );
    nor g1484 ( n1417 , n164 , n1435 );
    or g1485 ( n1724 , n1427 , n494 );
    xnor g1486 ( n1118 , n1086 , n842 );
    xnor g1487 ( n612 , n1037 , n848 );
    or g1488 ( n1063 , n490 , n1061 );
    or g1489 ( n1524 , n1316 , n607 );
    xnor g1490 ( n1098 , n410 , n663 );
    or g1491 ( n1482 , n1715 , n338 );
    and g1492 ( n390 , n315 , n1248 );
    xnor g1493 ( n781 , n987 , n1622 );
    and g1494 ( n323 , n975 , n1574 );
    and g1495 ( n198 , n1643 , n1707 );
    and g1496 ( n1281 , n1024 , n709 );
    nor g1497 ( n740 , n353 , n1360 );
    not g1498 ( n1768 , n1642 );
    or g1499 ( n7 , n182 , n595 );
    or g1500 ( n963 , n371 , n266 );
    or g1501 ( n1611 , n1422 , n159 );
    not g1502 ( n18 , n1709 );
    xnor g1503 ( n1714 , n509 , n964 );
    not g1504 ( n1069 , n949 );
    not g1505 ( n104 , n407 );
    and g1506 ( n817 , n1242 , n7 );
    not g1507 ( n1479 , n303 );
    xnor g1508 ( n724 , n258 , n145 );
    xnor g1509 ( n730 , n564 , n1372 );
    or g1510 ( n987 , n1411 , n1572 );
    nor g1511 ( n445 , n1722 , n772 );
    xnor g1512 ( n1347 , n993 , n1753 );
    or g1513 ( n945 , n1107 , n822 );
    and g1514 ( n326 , n586 , n136 );
    and g1515 ( n375 , n1554 , n124 );
    xnor g1516 ( n1750 , n180 , n622 );
    xnor g1517 ( n1010 , n1443 , n444 );
    and g1518 ( n542 , n1251 , n1345 );
    or g1519 ( n295 , n0 , n1618 );
    not g1520 ( n646 , n1155 );
    xnor g1521 ( n438 , n1607 , n931 );
    not g1522 ( n1089 , n927 );
    not g1523 ( n780 , n1376 );
    xnor g1524 ( n203 , n1107 , n700 );
    not g1525 ( n1193 , n736 );
    nor g1526 ( n80 , n1423 , n1316 );
    not g1527 ( n1593 , n1060 );
    or g1528 ( n1453 , n140 , n553 );
    or g1529 ( n214 , n739 , n734 );
    nor g1530 ( n640 , n1381 , n1006 );
    not g1531 ( n250 , n1541 );
    not g1532 ( n1072 , n1757 );
    and g1533 ( n283 , n369 , n733 );
    and g1534 ( n82 , n1057 , n463 );
    or g1535 ( n1566 , n1229 , n1591 );
    and g1536 ( n1540 , n155 , n266 );
    not g1537 ( n1361 , n1459 );
    xnor g1538 ( n407 , n501 , n708 );
    not g1539 ( n515 , n1033 );
    xnor g1540 ( n1120 , n996 , n1051 );
    nor g1541 ( n1291 , n154 , n970 );
    and g1542 ( n745 , n949 , n1071 );
    not g1543 ( n1255 , n647 );
    nor g1544 ( n1092 , n1659 , n1197 );
    and g1545 ( n1389 , n1754 , n25 );
    xnor g1546 ( n1578 , n934 , n732 );
    xnor g1547 ( n989 , n1137 , n1299 );
    and g1548 ( n1225 , n649 , n1182 );
    not g1549 ( n1726 , n1039 );
    or g1550 ( n758 , n266 , n887 );
    nor g1551 ( n554 , n1252 , n418 );
    not g1552 ( n342 , n1297 );
    or g1553 ( n628 , n127 , n1298 );
    xnor g1554 ( n319 , n805 , n764 );
    and g1555 ( n149 , n439 , n1320 );
    not g1556 ( n61 , n1009 );
    or g1557 ( n1254 , n1607 , n576 );
    xnor g1558 ( n944 , n1042 , n904 );
    or g1559 ( n1533 , n763 , n841 );
    xnor g1560 ( n1584 , n1448 , n1360 );
    and g1561 ( n1094 , n1447 , n940 );
    or g1562 ( n1097 , n746 , n1031 );
    not g1563 ( n1520 , n827 );
    and g1564 ( n147 , n1461 , n266 );
    and g1565 ( n425 , n901 , n992 );
    not g1566 ( n1426 , n547 );
    nor g1567 ( n1293 , n971 , n1396 );
    xnor g1568 ( n1151 , n1468 , n1445 );
    xnor g1569 ( n263 , n584 , n516 );
    nor g1570 ( n102 , n353 , n498 );
    not g1571 ( n587 , n1424 );
    or g1572 ( n1483 , n937 , n917 );
    not g1573 ( n798 , n745 );
    or g1574 ( n11 , n835 , n153 );
    not g1575 ( n230 , n706 );
    not g1576 ( n1663 , n1619 );
    or g1577 ( n1616 , n46 , n940 );
    or g1578 ( n672 , n1381 , n621 );
    xnor g1579 ( n248 , n353 , n1351 );
    or g1580 ( n412 , n777 , n186 );
    xnor g1581 ( n700 , n952 , n414 );
    not g1582 ( n1034 , n1751 );
    or g1583 ( n1370 , n666 , n365 );
    and g1584 ( n1114 , n1230 , n4 );
    xnor g1585 ( n1734 , n12 , n1176 );
    and g1586 ( n1362 , n1582 , n72 );
    not g1587 ( n667 , n347 );
    or g1588 ( n226 , n809 , n1732 );
    not g1589 ( n1183 , n1237 );
    or g1590 ( n1261 , n825 , n1164 );
    not g1591 ( n1661 , n531 );
    or g1592 ( n1674 , n1532 , n1641 );
    nor g1593 ( n866 , n26 , n296 );
    not g1594 ( n413 , n307 );
    and g1595 ( n768 , n1422 , n1624 );
    or g1596 ( n431 , n1488 , n1011 );
    not g1597 ( n394 , n318 );
    not g1598 ( n926 , n1263 );
    xnor g1599 ( n785 , n555 , n788 );
    or g1600 ( n1732 , n1072 , n487 );
    not g1601 ( n629 , n681 );
    and g1602 ( n1440 , n643 , n990 );
    or g1603 ( n512 , n1604 , n818 );
    or g1604 ( n466 , n1468 , n1700 );
    and g1605 ( n847 , n807 , n1439 );
    not g1606 ( n362 , n1655 );
    xnor g1607 ( n510 , n1546 , n263 );
    xnor g1608 ( n269 , n544 , n1642 );
    not g1609 ( n416 , n179 );
    nor g1610 ( n1695 , n165 , n1354 );
    nor g1611 ( n1035 , n870 , n402 );
    nor g1612 ( n705 , n837 , n1143 );
    xnor g1613 ( n1579 , n272 , n857 );
    xnor g1614 ( n689 , n1604 , n716 );
    or g1615 ( n264 , n720 , n518 );
    and g1616 ( n1617 , n247 , n201 );
    or g1617 ( n205 , n203 , n1270 );
    xnor g1618 ( n891 , n1165 , n707 );
    or g1619 ( n1583 , n143 , n1285 );
    xnor g1620 ( n103 , n1280 , n787 );
    nor g1621 ( n363 , n1219 , n1672 );
    nor g1622 ( n52 , n1770 , n4 );
    nor g1623 ( n1627 , n1329 , n1000 );
    or g1624 ( n797 , n1558 , n1212 );
    or g1625 ( n998 , n363 , n1309 );
    and g1626 ( n635 , n62 , n598 );
    xor g1627 ( n106 , n156 , n95 );
    not g1628 ( n1598 , n1672 );
    not g1629 ( n773 , n1543 );
    or g1630 ( n709 , n1527 , n1616 );
    xnor g1631 ( n575 , n1280 , n1217 );
    and g1632 ( n311 , n1765 , n502 );
    xnor g1633 ( n1393 , n1656 , n1064 );
    xor g1634 ( n1472 , n335 , n557 );
    or g1635 ( n1038 , n1761 , n313 );
    and g1636 ( n854 , n613 , n679 );
    nor g1637 ( n415 , n952 , n1296 );
    nor g1638 ( n1355 , n1422 , n266 );
    or g1639 ( n1019 , n108 , n1419 );
    or g1640 ( n1547 , n1504 , n434 );
    xnor g1641 ( n1032 , n562 , n1578 );
    xnor g1642 ( n602 , n111 , n1136 );
    xor g1643 ( n126 , n580 , n1385 );
    or g1644 ( n176 , n1000 , n690 );
    and g1645 ( n1427 , n1735 , n85 );
    xnor g1646 ( n613 , n1493 , n1747 );
    nor g1647 ( n913 , n1513 , n1167 );
    not g1648 ( n1564 , n749 );
    not g1649 ( n663 , n993 );
    xnor g1650 ( n949 , n1607 , n684 );
    and g1651 ( n692 , n1223 , n250 );
    or g1652 ( n1465 , n1059 , n818 );
    xnor g1653 ( n1262 , n1576 , n24 );
    nor g1654 ( n1358 , n1174 , n351 );
    or g1655 ( n1036 , n1428 , n1125 );
    not g1656 ( n845 , n1364 );
    not g1657 ( n1612 , n1717 );
    or g1658 ( n922 , n359 , n327 );
    or g1659 ( n1412 , n520 , n1210 );
    or g1660 ( n1551 , n266 , n1648 );
    not g1661 ( n132 , n1253 );
    not g1662 ( n64 , n93 );
    or g1663 ( n860 , n681 , n1560 );
    or g1664 ( n1313 , n530 , n377 );
    and g1665 ( n974 , n35 , n907 );
    xnor g1666 ( n1752 , n914 , n138 );
    xnor g1667 ( n1525 , n1719 , n1683 );
    not g1668 ( n1153 , n1296 );
    not g1669 ( n1160 , n585 );
    not g1670 ( n196 , n1075 );
    xnor g1671 ( n1204 , n666 , n288 );
    xnor g1672 ( n40 , n210 , n17 );
    xnor g1673 ( n670 , n816 , n138 );
    or g1674 ( n420 , n1000 , n1281 );
    xnor g1675 ( n1717 , n1744 , n1459 );
    not g1676 ( n516 , n386 );
    buf g1677 ( n292 , n1677 );
    or g1678 ( n1478 , n377 , n1167 );
    nor g1679 ( n110 , n353 , n98 );
    not g1680 ( n145 , n428 );
endmodule
